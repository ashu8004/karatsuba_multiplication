module partial_products(input  [15:0]a,input  [15:0]b,output reg [31:0]p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
always @(a or b)
	begin
		p0<=b[0]?a:32'b0;
		p1<=b[1]?(a<<1):32'b0;
		p2<=b[2]?(a<<2):32'b0;
		p3<=b[3]?(a<<3):32'b0;
		p4<=b[4]?(a<<4):32'b0;
		p5<=b[5]?(a<<5):32'b0;
		p6<=b[6]?(a<<6):32'b0;
		p7<=b[7]?(a<<7):32'b0;
		p8<=b[8]?(a<<8):32'b0;
		p9<=b[9]?(a<<9):32'b0;
		p10<=b[10]?(a<<10):32'b0;
		p11<=b[11]?(a<<11):32'b0;
		p12<=b[12]?(a<<12):32'b0;
		p13<=b[13]?(a<<13):32'b0;
		p14<=b[14]?(a<<14):32'b0;
		p15<=b[15]?(a<<15):32'b0;
	end
endmodule
